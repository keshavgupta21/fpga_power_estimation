module top(
    input wire clk100mhz,
    output wire [3:0] led
);

endmodule