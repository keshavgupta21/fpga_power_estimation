module user(
    input wire clk100m,
    input wire rstn
);

endmodule