module top(
    input wire clk100m,
    output wire [3:0] led
);

endmodule